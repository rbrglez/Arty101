---------------------------------------------------------------------------------------------------
--! @brief
--!
--! @author
--!
--! @date 
--!
--! @version v0.1
--!
--! @file MarkDebugPkg.vhd
--!
---------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;
library surf;
use surf.StdRtlPkg.all;

package MarkDebugPkg is

   -- Marked for debug
   constant TOP_DEBUG_C : string := "false";

end MarkDebugPkg;

package body MarkDebugPkg is
end MarkDebugPkg;
