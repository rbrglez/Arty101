----------------------------------------------------------------------------------------------------
-- @brief VgaDisplayArtyTestPkg
--
-- @author Rene Brglez (rene.brglez@gmail.com)
--
-- @date December 2022
-- 
-- @version v0.1
--
-- @file VgaDisplayArtyTestPkg.vhd
--
----------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;
library surf;
use surf.StdRtlPkg.all;

package VgaDisplayArtyTestPkg is

   constant CLK_FREQ_C : real := 100.0E6;

end VgaDisplayArtyTestPkg;

package body VgaDisplayArtyTestPkg is

end package body VgaDisplayArtyTestPkg;
