----------------------------------------------------------------------------------------------------
-- @brief SegmentDisplayArtyTestPkg
--
-- @author Rene Brglez (rene.brglez@gmail.com)
--
-- @date December 2022
-- 
-- @version v0.1
--
-- @file SegmentDisplayArtyTestPkg.vhd
--
----------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;
use work.StdRtlPkg.all;

package SegmentDisplayArtyTestPkg is

end SegmentDisplayArtyTestPkg;

package body SegmentDisplayArtyTestPkg is

end package body SegmentDisplayArtyTestPkg;
