----------------------------------------------------------------------------------------------------
-- @brief ArtySegmentDisplayTestPkg
--
-- @author Rene Brglez (rene.brglez@gmail.com)
--
-- @date December 2022
-- 
-- @version v0.1
--
-- @file ArtySegmentDisplayTestPkg.vhd
--
----------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;
library surf;
use surf.StdRtlPkg.all;

package ArtySegmentDisplayTestPkg is

   constant CLK_FREQ_C : real := 100.0E6;

end ArtySegmentDisplayTestPkg;

package body ArtySegmentDisplayTestPkg is

end package body ArtySegmentDisplayTestPkg;
